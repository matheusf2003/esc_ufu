module add16(input [15:0] a, input [15:0] b, output [0:15] sum);
    assign sum = a + b;

endmodule