//
// Multiplexador de duas entradas (16 bits), comportamental
//
module mux4way16(input [15:0] a, input [15:0] b, input [15:0] c, input [15:0] d, input [1:0] sel, output [15:0] y);

  assign y = (sel == 2'b00) ? a :
    (sel == 2'b01) ? b :
    (sel == 2'b10) ? c : d;

endmodule

